`timescale 1us/1ns

module 
